----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/28/2023 01:04:20 AM
-- Design Name: 
-- Module Name: coef - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity coef is
    Port ( clk : in std_logic;
           segment : in STD_LOGIC_VECTOR (7 downto 0);
           c0 : out unsigned (18 downto 0);
           c1 : out signed (17 downto 0);
           c2 : out unsigned (17 downto 0));
end coef;

architecture Behavioral of coef is
signal data : unsigned (54 downto 0);

begin

proc_sense: process(segment)
begin
    case segment is
        when "00000000" => data <= "0000010101100101001100110111110001110010100011110000000";
        when "00000001" => data <= "0000001111101000111101001011111011001001011111011110011";
        when "00000010" => data <= "0000001010001100100101010111101101110000110010101000000";
        when "00000011" => data <= "0000000101000010001101011101111111001000001111111010011";
        when "00000100" => data <= "0000100100110011110101100101100100010010101101110011100";
        when "00000101" => data <= "0000100000010100011101111010111110111001110101000001100";
        when "00000110" => data <= "0000011100011000111110001001011101011001010011011010011";
        when "00000111" => data <= "0000011000110110001110010011110011100000111101101011001";
        when "00001000" => data <= "0000110001000101110101111110110101010010100011001000110";
        when "00001001" => data <= "0000101101010111101110010010111100001001101111010111011";
        when "00001010" => data <= "0000101010001011010110100000101110001001010000111111000";
        when "00001011" => data <= "0000100111010110110110101010110001001000111101100100011";
        when "00001100" => data <= "0000111011100110110110001111001100101010010111001100011";
        when "00001101" => data <= "0000111000010111111110100001110101001001100111010010101";
        when "00001110" => data <= "0000110101101000010110101110100111010001001011010000101";
        when "00001111" => data <= "0000110011001110111110110111111100110000111001011001010";
        when "00010000" => data <= "0001000100111011000110011010110100101010001100100110110";
        when "00010001" => data <= "0001000010000010000110101100001001100001011111111010010";
        when "00010010" => data <= "0000111111100110010110111000000001000001000101110011111";
        when "00010011" => data <= "0000111101011110111111000000101011011000110101001101001";
        when "00010100" => data <= "0001001101010111000110100011100101111010000011100100011";
        when "00010101" => data <= "0001001010101110100110110011110011100001011001100101001";
        when "00010110" => data <= "0001001000100001010110111110111000110001000001000110100";
        when "00010111" => data <= "0001000110100111000111000110111101101000110001100011100";
        when "00011000" => data <= "0001010101000111110110101010011111110001111011110111110";
        when "00011001" => data <= "0001010010101100000110111001110000100001010100001100011";
        when "00011010" => data <= "0001010000101010000111000100001011001000111101000110010";
        when "00011011" => data <= "0001001110111001111111001011110000001000101110011100100";
        when "00011100" => data <= "0001011100010101101110110000000110101001110101010001000";
        when "00011101" => data <= "0001011010000100011110111110100011001001001111100101010";
        when "00011110" => data <= "0001011000001011011111001000011001010000111001101011010";
        when "00011111" => data <= "0001010110100011010111001111100011001000101011110010110";
        when "00100000" => data <= "0001100011000111001110110100110001001001101111100010101";
        when "00100001" => data <= "0001100000111110011111000010100000101001001011100110010";
        when "00100010" => data <= "0001011111001100110111001011110111001000110110101110100";
        when "00100011" => data <= "0001011101101011011111010010101001100000101001100000110";
        when "00100100" => data <= "0001101001100000100110111000101110100001101010100010001";
        when "00100101" => data <= "0001100111011111001111000101110110010001001000000111110";
        when "00100110" => data <= "0001100101110011110111001110110001010000110100001010001";
        when "00100111" => data <= "0001100100010111110111010101001111011000100111100001111";
        when "00101000" => data <= "0001101111100101100110111100001000101001100110000110111";
        when "00101001" => data <= "0001101101101010011111001000101101101001000101000011110";
        when "00101010" => data <= "0001101100000100011111010001010000011000110001111001101";
        when "00101011" => data <= "0001101010101101000111010111011100011000100101110010101";
        when "00101100" => data <= "0001110101011000101110111111000111001001100010001010110";
        when "00101101" => data <= "0001110011100011000111001011001101000001000010010101101";
        when "00101110" => data <= "0001110010000001101111010011011010001000101111111001101";
        when "00101111" => data <= "0001110000101110011111011001010110011000100100010000001";
        when "00110000" => data <= "0001111010111100001111000001101111010001011110101000100";
        when "00110001" => data <= "0001111001001011011111001101011001001000111111111001110";
        when "00110010" => data <= "0001110111101110000111010101010011000000101110000111001";
        when "00110011" => data <= "0001110110011110011111011011000001000000100010111000010";
        when "00110100" => data <= "0010000000010001111111000100000100111001011011011100010";
        when "00110101" => data <= "0001111110100101011111001111010101101000111101101101001";
        when "00110110" => data <= "0001111101001011101111010110111110001000101100100000001";
        when "00110111" => data <= "0001111011111111001111011100011111010000100001101001010";
        when "00111000" => data <= "0010000101011011010111000110001011010001011000100010101";
        when "00111001" => data <= "0010000011110010100111010001000101001000111011101101101";
        when "00111010" => data <= "0010000010011100000111011000011101110000101011000010110";
        when "00111011" => data <= "0010000001010010010111011101110011011000100000100001110";
        when "00111100" => data <= "0010001010011001011111001000000100110001010101111001000";
        when "00111101" => data <= "0010001000110100001111010010101001110000111001111001011";
        when "00111110" => data <= "0010000111100000101111011001110100000000101001101101110";
        when "00111111" => data <= "0010000110011001011111011110111111001000011111100000110";
        when "01000000" => data <= "0010001111001101011111001001110011010001010011011101011";
        when "01000001" => data <= "0010001101101011010111010100000101000000111000001110110";
        when "01000010" => data <= "0010001100011010011111011011000010001000101000011111111";
        when "01000011" => data <= "0010001011010101100111100000000011100000011110100101010";
        when "01000100" => data <= "0010010011111000010111001011011000010001010001001101111";
        when "01000101" => data <= "0010010010011001000111010101011000011000110110101100101";
        when "01000110" => data <= "0010010001001010100111011100001001011000100111011000011";
        when "01000111" => data <= "0010010000000111110111100001000001111000011101101110101";
        when "01001000" => data <= "0010011000011010100111001100110101010001001111001001001";
        when "01001001" => data <= "0010010110111110000111010110100101000000110101010001111";
        when "01001010" => data <= "0010010101110001110111011101001010101000100110010110010";
        when "01001011" => data <= "0010010100110000111111100001111011000000011100111100001";
        when "01001100" => data <= "0010011100110101001111001110001011000001001101001101110";
        when "01001101" => data <= "0010011011011011000111010111101011100000110011111101110";
        when "01001110" => data <= "0010011010010000110111011110000110110000100101011000111";
        when "01001111" => data <= "0010011001010001101111100010101111100000011100001101100";
        when "01010000" => data <= "0010100001001000100111001111011010100001001011011010110";
        when "01010001" => data <= "0010011111110000101111011000101100111000110010101111010";
        when "01010010" => data <= "0010011110101000010111011110111110011000100100011111111";
        when "01010011" => data <= "0010011101101010110111100011100000001000011011100010000";
        when "01010100" => data <= "0010100101010101001111010000100100011001001001101111010";
        when "01010101" => data <= "0010100011111111011111011001101001100000110001100110000";
        when "01010110" => data <= "0010100010111000110111011111110010000000100011101010101";
        when "01010111" => data <= "0010100001111100110111100100001101001000011010111001100";
        when "01011000" => data <= "0010101001011011100111010001101001011001001000001010100";
        when "01011001" => data <= "0010101000000111110111011010100010000000110000100001100";
        when "01011010" => data <= "0010100111000010110111100000100010001000100010111000110";
        when "01011011" => data <= "0010100110001000001111100100110111000000011010010011100";
        when "01011100" => data <= "0010101101011100000111010010101001111001000110101011110";
        when "01011101" => data <= "0010101100001010001111011011010111000000101111100001000";
        when "01011110" => data <= "0010101011000110110111100001001111000000100010001010000";
        when "01011111" => data <= "0010101010001101011111100101011110001000011001110000000";
        when "01100000" => data <= "0010110001010111001111010011100110100001000101010010101";
        when "01100001" => data <= "0010110000000110111111011100001000100000101110100100011";
        when "01100010" => data <= "0010101111000101000111100001111001001000100001011110000";
        when "01100011" => data <= "0010101110001100111111100110000010110000011001001110100";
        when "01100100" => data <= "0010110101001101001111010100011111100001000011111110011";
        when "01100101" => data <= "0010110011111110100111011100110111001000101101101011001";
        when "01100110" => data <= "0010110010111101111111100010100000101000100000110100100";
        when "01100111" => data <= "0010110010000111000111100110100101001000011000101111000";
        when "01101000" => data <= "0010111000111110010111010101010101010001000010101110101";
        when "01101001" => data <= "0010110111110001010111011101100011001000101100110101000";
        when "01101010" => data <= "0010110110110001111111100011000101111000100000001101010";
        when "01101011" => data <= "0010110101111100000111100111000101100000011000010001010";
        when "01101100" => data <= "0010111100101010111111010110001000000001000001100011001";
        when "01101101" => data <= "0010111011011111010111011110001100101000101100000001110";
        when "01101110" => data <= "0010111010100001000111100011101001000000011111101000001";
        when "01101111" => data <= "0010111001101100010111100111100100000000010111110101000";
        when "01110000" => data <= "0011000000010011001111010110111000001001000000011011011";
        when "01110001" => data <= "0010111111001000111111011110110011111000101011010001001";
        when "01110010" => data <= "0010111110001011110111100100001010011000011111000100111";
        when "01110011" => data <= "0010111101011000000111101000000000111000010111011010010";
        when "01110100" => data <= "0011000011110111010111010111100101110000111111010111001";
        when "01110101" => data <= "0011000010101110010111011111011001001000101010100010111";
        when "01110110" => data <= "0011000001110010011111100100101001111000011110100011011";
        when "01110111" => data <= "0011000000111111011111101000011100010000010111000000111";
        when "01111000" => data <= "0011000111010111100111011000010001010000111110010110001";
        when "01111001" => data <= "0011000110001111110111011111111100100000101001110110111";
        when "01111010" => data <= "0011000101010100111111100101000111110000011110000011100";
        when "01111011" => data <= "0011000100100010110111101000110110010000010110101000110";
        when "01111100" => data <= "0011001010110100001111011000111010100000111101011000001";
        when "01111101" => data <= "0011001001101101100111100000011110001000101001001100110";
        when "01111110" => data <= "0011001000110011100111100101100100010000011101100101001";
        when "01111111" => data <= "0011001000000010011111101001001111000000010110010001110";
        when "10000000" => data <= "0011001110001101001111011001100001111000111100011100111";
        when "10000001" => data <= "0011001101000111101111100000111110010000101000100100101";
        when "10000010" => data <= "0011001100001110101111100101111111011000011101001000001";
        when "10000011" => data <= "0011001011011110010111101001100110100000010101111011110";
        when "10000100" => data <= "0011010001100010110111011010000111100000111011100100001";
        when "10000101" => data <= "0011010000011110011111100001011100111000100111111110010";
        when "10000110" => data <= "0011001111100110010111100110011001001000011100101100011";
        when "10000111" => data <= "0011001110110110101111101001111100111000010101100110101";
        when "10001000" => data <= "0011010100110101010111011010101011011000111010101101111";
        when "10001001" => data <= "0011010011110001111111100001111010001000100111011001101";
        when "10001010" => data <= "0011010010111010101111100110110001111000011100010001111";
        when "10001011" => data <= "0011010010001011101111101010010010010000010101010010101";
        when "10001100" => data <= "0011011000000100101111011011001101110000111001111001110";
        when "10001101" => data <= "0011010111000010010111100010010110001000100110110110011";
        when "10001110" => data <= "0011010110001011110111100111001001100000011011111000011";
        when "10001111" => data <= "0011010101011101100111101010100110110000010100111111010";
        when "10010000" => data <= "0011011011010001001111011011101110110000111001000111110";
        when "10010001" => data <= "0011011010001111101111100010110000111000100110010100100";
        when "10010010" => data <= "0011011001011001111111100111100000001000011011100000000";
        when "10010011" => data <= "0011011000101100010111101010111010011000010100101100111";
        when "10010100" => data <= "0011011110011010110111011100001110011000111000010111101";
        when "10010101" => data <= "0011011101011010001111100011001010101000100101110100000";
        when "10010110" => data <= "0011011100100101001111100111110101111000011011001000100";
        when "10010111" => data <= "0011011011111000010111101011001101010000010100011011000";
        when "10011000" => data <= "0011100001100001101111011100101100111000110111101001100";
        when "10011001" => data <= "0011100000100001111111100011100011011000100101010100110";
        when "10011010" => data <= "0011011111101101101111101000001010110000011010110001111";
        when "10011011" => data <= "0011011111000001010111101011011111010000010100001010000";
        when "10011100" => data <= "0011100100100110000111011101001010001000110110111100111";
        when "10011101" => data <= "0011100011100111000111100011111011001000100100110110110";
        when "10011110" => data <= "0011100010110011100111101000011110110000011010011100010";
        when "10011111" => data <= "0011100010000111110111101011110000101000010011111001101";
        when "10100000" => data <= "0011100111100111110111011101100110010000110110010010000";
        when "10100001" => data <= "0011100110101001101111100100010001111000100100011001110";
        when "10100010" => data <= "0011100101110110110111101000110010000000011010000111010";
        when "10100011" => data <= "0011100101001011100111101100000001010000010011101001110";
        when "10100100" => data <= "0011101010100111001111011110000001011000110101101000101";
        when "10100101" => data <= "0011101001101001110111100100101000000000100011111101110";
        when "10100110" => data <= "0011101000110111100111101001000100101000011001110011001";
        when "10100111" => data <= "0011101000001100111111101100010001010000010011011010100";
        when "10101000" => data <= "0011101101100100001111011110011011100000110101000000101";
        when "10101001" => data <= "0011101100100111101111100100111101001000100011100010111";
        when "10101010" => data <= "0011101011110101111111101001010110100000011001011111101";
        when "10101011" => data <= "0011101011001011110111101100100000110000010011001011110";
        when "10101100" => data <= "0011110000011111000111011110110100110000110100011010000";
        when "10101101" => data <= "0011101111100011001111100101010001101000100011001000110";
        when "10101110" => data <= "0011101110110010000111101001100111110000011001001100111";
        when "10101111" => data <= "0011101110001000011111101100101111110000010010111101101";
        when "10110000" => data <= "0011110011010111101111011111001101001000110011110100110";
        when "10110001" => data <= "0011110010011100100111100101100101011000100010101111100";
        when "10110010" => data <= "0011110001101011111111101001111000011000011000111010110";
        when "10110011" => data <= "0011110001000010110111101100111110001000010010101111111";
        when "10110100" => data <= "0011110110001110001111011111100100101000110011010000101";
        when "10110101" => data <= "0011110101010011101111100101111000100000100010010111001";
        when "10110110" => data <= "0011110100100011101111101010001000100000011000101001001";
        when "10110111" => data <= "0011110011111011000111101101001100000000010010100010100";
        when "10111000" => data <= "0011111001000010110111011111111011011000110010101101101";
        when "10111001" => data <= "0011111000001000111111100110001011000000100001111111101";
        when "10111010" => data <= "0011110111011001011111101010011000000000011000011000001";
        when "10111011" => data <= "0011110110110001001111101101011001100000010010010101110";
        when "10111100" => data <= "0011111011110101010111100000010001100000110010001011110";
        when "10111101" => data <= "0011111010111100000111100110011100111000100001101000110";
        when "10111110" => data <= "0011111010001101001111101010100111001000011000000111101";
        when "10111111" => data <= "0011111001100101010111101101100110100000010010001001010";
        when "11000000" => data <= "0011111110100101111111100000100110111000110001101011000";
        when "11000001" => data <= "0011111101101101010111100110101110010000100001010010101";
        when "11000010" => data <= "0011111100111110111111101010110101101000010111110111110";
        when "11000011" => data <= "0011111100010111100111101101110011001000010001111101010";
        when "11000100" => data <= "0100000001010100110111100000111011101000110001001011010";
        when "11000101" => data <= "0100000000011100101111100110111111000000100000111101010";
        when "11000110" => data <= "0011111111101110110111101011000011110000010111101000010";
        when "11000111" => data <= "0011111111000111110111101101111111010000010001110001100";
        when "11001000" => data <= "0100000100000001110111100001001111101000110000101100101";
        when "11001001" => data <= "0100000011001010010111100111001111010000100000101000100";
        when "11001010" => data <= "0100000010011100110111101011010001100000010111011001011";
        when "11001011" => data <= "0100000001110110010111101110001011001000010001100110010";
        when "11001100" => data <= "0100000110101101001111100001100011001000110000001111001";
        when "11001101" => data <= "0100000101110110001111100111011111000000100000010100101";
        when "11001110" => data <= "0100000101001001001111101011011110110000010111001011000";
        when "11001111" => data <= "0100000100100011000111101110010110101000010001011011011";
        when "11010000" => data <= "0100001001010110110111100001110110000000101111110011010";
        when "11010001" => data <= "0100001000100000010111100111101110011000100000000001101";
        when "11010010" => data <= "0100000111110011110111101011101011101000010110111101010";
        when "11010011" => data <= "0100000111001101111111101110100001110000010001010001000";
        when "11010100" => data <= "0100001011111110110111100010001000010000101111011001100";
        when "11010101" => data <= "0100001011001000111111100111111101001000011111101111111";
        when "11010110" => data <= "0100001010011100101111101011111000001000010110110000010";
        when "11010111" => data <= "0100001001110111010111101110101100100000010001000111001";
        when "11011000" => data <= "0100001110100101001111100010011001110000101111000011000";
        when "11011001" => data <= "0100001101101111110111101000001011100000011111100000001";
        when "11011010" => data <= "0100001101000100000111101100000100010000010110100100101";
        when "11011011" => data <= "0100001100011110111111101110110111000000010000111110001";
        when "11011100" => data <= "0100010001001010000111100010101010100000101110110010010";
        when "11011101" => data <= "0100010000010101001111101000011001010000011111010011101";
        when "11011110" => data <= "0100001111101001110111101100001111111000010110011011000";
        when "11011111" => data <= "0100001111000101000111101111000001001000010000110110100";
        when "11100000" => data <= "0100010011101101011111100010111010010000101110101100100";
        when "11100001" => data <= "0100010010111000111111101000100110010000011111001101001";
        when "11100010" => data <= "0100010010001110000111101100011011000000010110010101000";
        when "11100011" => data <= "0100010001101001101111101111001010110000010000110001010";
        when "11100100" => data <= "0100010110001111010111100011001000101000101110111011101";
        when "11100101" => data <= "0100010101011011010111101000110010011000011111010010001";
        when "11100110" => data <= "0100010100110000110111101100100101100000010110010110000";
        when "11100111" => data <= "0100010100001100101111101111010100000000010000110000101";
        when "11101000" => data <= "0100011000101111110111100011010100111000101111110100001";
        when "11101001" => data <= "0100010111111100010111101000111101011000011111101101110";
        when "11101010" => data <= "0100010111010010000111101100101111001000010110100100111";
        when "11101011" => data <= "0100010110101110010111101111011100101000010000111001000";
        when "11101100" => data <= "0100011011001110111111100101000100000000000000000000000";
        when "11101101" => data <= "0100011010011011110111101010001001010000000000000000000";
        when "11101110" => data <= "0100011001110010000111101101100110110000000000000000000";
        when "11101111" => data <= "0100011001001110100111110000000111011000000000000000000";
        when "11110000" => data <= "0100011101101100101000000000000000000000000000000000000";
        when "11110001" => data <= "0100011100111010000000000000000000000000000000000000000";
        when "11110010" => data <= "0100011100010000100000000000000000000000000000000000000";
        when "11110011" => data <= "0100011011101101011000000000000000000000000000000000000";
        when "11110100" => data <= "0100100100111110000000000000000000000000000000000000000";
        when "11110101" => data <= "0100100010100100001000000000000000000000000000000000000";
        when "11110110" => data <= "0100100000001001000000000000000000000000000000000000000";
        when "11110111" => data <= "0100011110101101101000000000000000000000000000000000000";
        when others => data <= "0000000000000000000000000000000000000000000000000000000";
    end case; 
end process proc_sense;

proc_dataout: process(clk)
begin
    if rising_edge(clk) then
            c0 <= data(54 downto 36);
            c1 <= signed(data(35 downto 18));
            c2 <= data(17 downto 0);
    end if;
end process proc_dataout;

end Behavioral;
